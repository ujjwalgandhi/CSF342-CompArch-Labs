module magcomp(out, a, b);
	input [3:0]a, [3:0]b;
	output [1:0] c;
	
endmodule